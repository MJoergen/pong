library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
    
package sprite_pkg is
    type pattern_t is array (integer range 0 to 20) of std_logic_vector(0 to 23);
end package sprite_pkg;

